Require Import ssreflect ssrbool ssrfun eqtype fintype finfun finset ssralg.
Require Import bigop seq choice ssrnat prime ssralg fingroup pgroup zmodp.
Require Import matrix vector galgebra algebra.

(*****************************************************************************)
(*  * Module over an algebra                                                 *)
(*     amoduleType A    == type for finite dimension module structure.       *)
(*                                                                           *)
(*        v :* x        == right product of the module                       *)
(*      (M :* A)%VS     == the smallest vector space that contains           *)
(*                           {v :* x | v \in M & x \in A}                    *)
(*      (modv M A)      == M is a module for A                               *)
(*      (modf f M A)    == f is a module homomorphism on M for A             *)
(*****************************************************************************)
(*****************************************************************************)

Set Implicit Arguments.
Unset Strict Implicit.
Unset Printing Implicit Defensive.
Open Local Scope ring_scope.

Delimit Scope amodule_scope with aMS.

Import GRing.Theory.

Module AModuleType.
Section ClassDef.

Variable R : ringType.
Variable V: vspaceType R.
Variable A: algFType R.

Structure mixin_of (V : vspaceType R) : Type := Mixin {
  action: A -> 'End(V);
  action_morph: forall x a b, action (a * b) x = action b (action a x);
  action_linear: forall x , linear (action^~ x);
  action1: forall x , action 1 x = x 
}.

Structure class_of (V : Type) : Type := Class {
  base : VectorType.class_of R V;
   mixin : mixin_of (VectorType.Pack _ base V) 
}.
Local Coercion base : class_of >-> VectorType.class_of.

Implicit Type phA : phant A.

Structure type phA : Type := Pack {sort : Type; _ : class_of sort; _ : Type}.
Local Coercion sort : type >-> Sortclass.

Definition class phA (cT : type phA):=
  let: Pack _ c _ := cT return class_of cT in c.
Definition clone phA T cT c of phant_id (@class phA cT) c := @Pack phA T c T.

Definition pack phA V V0 (m0 : mixin_of (@VectorType.Pack R _ V V0 V)) :=
  fun bT b & phant_id (@VectorType.class _ (Phant R) bT) b =>
  fun    m & phant_id m0 m => Pack phA (@Class V b m) V.

Definition eqType phA cT := Equality.Pack (@class phA cT) cT.
Definition choiceType phA cT := choice.Choice.Pack (@class phA cT) cT.
Definition zmodType phA cT := GRing.Zmodule.Pack (@class phA cT) cT.
Definition lmodType phA cT := GRing.Lmodule.Pack (Phant R) (@class phA cT) cT.
Definition vectType phA cT := VectorType.Pack (Phant R) (@class phA cT) cT.

End ClassDef.

Module Exports.
Coercion base : class_of >->  VectorType.class_of.
Coercion mixin : class_of >-> mixin_of.
Coercion sort : type >-> Sortclass.

Coercion eqType : type >->  Equality.type.
Canonical Structure eqType.
Coercion choiceType : type >-> Choice.type.
Canonical Structure choiceType.
Coercion zmodType : type >-> GRing.Zmodule.type.
Canonical Structure zmodType.
Coercion lmodType : type>->  GRing.Lmodule.type.
Canonical Structure lmodType.
Coercion vectType : type >-> VectorType.type.
Canonical Structure vectType.

Notation amoduleType A := (@type _ _ (Phant A)).
Notation AModuleType A m := (@pack _ _ (Phant A) _ _ m _ _ id _ id).
Notation AModuleMixin := Mixin.

Bind Scope ring_scope with sort.
End Exports.

End AModuleType.
Import AModuleType.Exports.

Section AModuleDef.
Variables (F : fieldType) (A: algFType F) (M: amoduleType A).

Definition rmorph (a: A) := AModuleType.action (AModuleType.class M) a.
Definition rmul (a: M) (b: A) : M := rmorph b a.
Notation "a :* b" := (rmul a b): ring_scope.

Implicit Types x y: A.
Implicit Types v w: M.
Implicit Types c: F.

Lemma rmulD x: {morph (rmul^~ x): v1 v2 / v1 + v2}.
Proof. move=> *; exact: linearD. Qed.

Lemma rmul_linear_proof : forall  v, linear (rmul v).
Proof. by rewrite /rmul /rmorph; case: M => s [] b []. Qed.
Canonical Structure rmul_linear v := GRing.Linear (rmul_linear_proof v).

Lemma rmulA v x y: v :* (x * y) = (v :* x) :* y.
Proof. exact: AModuleType.action_morph. Qed.

Lemma rmulZ : forall c v x, (c *: v) :* x = c *: (v :* x).
Proof. move=> c v x; exact: linearZ. Qed.

Lemma rmul0 : left_zero 0 rmul.
Proof. move=> x; exact: linear0. Qed.

Lemma rmul1 : forall v , v :* 1 = v.
Proof. by rewrite /rmul /rmorph; case: M => s [] b []. Qed.

Lemma rmul_sum :  forall I r P (f : I -> M) x,
  \sum_(i <- r | P i) f i :* x = (\sum_(i <- r | P i) f i) :* x.
Proof.
by move=> I r P f x; rewrite -linear_sum.
Qed.

Implicit Types vs: {vspace M}.
Implicit Types ws: {vspace A}.

Definition eprodv vs ws := span (allpairs rmul (vbasis vs) (vbasis ws)).
Local Notation "A :* B" := (eprodv A B) : vspace_scope.

Lemma memv_eprod : forall vs ws a b , a \in vs -> b \in ws -> a :* b \in (vs :* ws)%VS.
Proof. 
move=> vs ws a b Ha Hb.
rewrite (coord_basis Ha) (coord_basis Hb).
rewrite linear_sum /=; apply: memv_sum => [] [j Hj] _.
rewrite -rmul_sum; apply: memv_sum => [] [i Hi] _ /=.
rewrite linearZ memvZl //= rmulZ memvZl //=.
apply: memv_span; apply/allpairsP; exists ((vbasis vs)`_i, (vbasis ws)`_j)=> //.
by rewrite !mem_nth /=.
Qed.

Lemma eprodvP : forall vs1 ws vs2,   reflect (forall a b, a \in vs1 -> b \in ws -> a :* b \in vs2)
          (vs1 :* ws <= vs2)%VS.
Proof.
move=> vs1 ws vs2; apply: (iffP idP).
  move=> Hs a b Ha Hb.
  by apply: subsetv_trans Hs; exact: memv_eprod.
move=> Ha; apply/subsetvP=> v.
move/coord_span->; apply: memv_sum => [] [i /= Hi] _.
apply: memvZl; move: (mem_nth 0 Hi); case/allpairsP=> p [I1 I2 ->].
by rewrite Ha // memv_basis.
Qed.

Lemma eprod0v: left_zero (0%:VS) eprodv.
Proof.
move=> vs; apply subsetv_anti; rewrite subset0v andbT.
apply/eprodvP=> a b; case/injvP=> k1 -> Hb.
by rewrite scaler0 rmul0 mem0v.
Qed.

Lemma eprodv0 : forall vs, (vs :* 0%:VS = 0%:VS)%VS.
Proof.
move=> vs; apply subsetv_anti; rewrite subset0v andbT.
apply/eprodvP=> a b Ha; case/injvP=> k1 ->.
by rewrite scaler0 linear0 mem0v.
Qed.

Lemma eprodv1 : forall vs, (vs :* 1%:VS = vs)%VS.
Proof.
case: (vbasis1 A)=> k [Hk He] /=.
move=> vs; apply subsetv_anti; apply/andP; split.
  apply/eprodvP=> a b Ha; case/injvP=> k1 ->.
  by rewrite linearZ /= rmul1 memvZl.
apply/subsetvP=> v Hv.
rewrite (coord_basis Hv); apply: memv_sum => [] [i Hi] _ /=.  
apply: memvZl.
rewrite -[_`_i]rmul1; apply: memv_eprod; last by apply: memv_inj.
by apply: memv_basis; apply: mem_nth.
Qed.

Lemma eprodv_monol : forall ws vs1 vs2, (vs1 <= vs2 -> vs1 :* ws <= vs2 :* ws)%VS.
Proof.
move=> ws vs1 vs2 Hvs; apply/eprodvP=> a b Ha Hb; apply: memv_eprod=> //.
by apply: subsetv_trans Hvs.
Qed.

Lemma eprodv_monor : forall vs ws1 ws2, (ws1 <= ws2 -> vs :* ws1 <= vs :* ws2)%VS.
Proof.
move=> vs ws1 ws2 Hvs; apply/eprodvP=> a b Ha Hb; apply: memv_eprod=> //.
by apply: subsetv_trans Hvs.
Qed.

Lemma eprodv_addl: left_distributive eprodv addv.
Proof.
move=> vs1 vs2 ws; apply subsetv_anti; apply/andP; split.
  apply/eprodvP=> a b;case/addv_memP=> v1 [v2 [Hv1 Hv2 ->]] Hb.
  by rewrite rmulD; apply: addv_mem; apply: memv_eprod.
apply/subsetvP=> v;  case/addv_memP=> v1 [v2 [Hv1 Hv2 ->]].
apply: memvD.
  move: v1 Hv1; apply/subsetvP; apply: eprodv_monol; exact: addvSl.
move: v2 Hv2; apply/subsetvP; apply: eprodv_monol; exact: addvSr.
Qed.

Lemma eprodv_sumr : forall vs ws1 ws2, (vs :* (ws1 + ws2) = vs :* ws1 + vs :* ws2)%VS.
Proof.
move=> vs ws1 ws2; apply subsetv_anti; apply/andP; split.
  apply/eprodvP=> a b Ha;case/addv_memP=> v1 [v2 [Hv1 Hv2 ->]].
  by rewrite linearD; apply: addv_mem; apply: memv_eprod.
apply/subsetvP=> v;  case/addv_memP=> v1 [v2 [Hv1 Hv2 ->]].
apply: memvD.
  move: v1 Hv1; apply/subsetvP; apply: eprodv_monor; exact: addvSl.
move: v2 Hv2; apply/subsetvP; apply: eprodv_monor; exact: addvSr.
Qed.

Definition modv (vs: {vspace M}) (al: {algebra A}) :=
   (vs :* al  <= vs)%VS.
 
Lemma mod0v : forall al , modv 0%:VS al.
Proof. by move=> al; rewrite /modv eprod0v subsetv_refl. Qed.

Lemma modv1 : forall vs , modv vs (aspace1 A).
Proof. by move=> vs; rewrite /modv eprodv1 subsetv_refl. Qed.

Lemma modfv : forall al,  modv (fullv M) al.
Proof. by move=> al; exact: subsetvf. Qed.

Lemma memv_mod_mul : forall ms al m a, 
  modv ms al -> m \in ms -> a \in al -> m :* a \in ms.
Proof. 
move=> ms al m a Hmo Hm Ha; apply: subsetv_trans Hmo.
by apply: memv_eprod.
Qed.

Lemma modvD : forall ms1 ms2 al , 
  modv ms1 al -> modv ms2 al -> modv (ms1 + ms2)%VS al.
Proof.
move=> ms1 ms2 al Hm1 Hm2; rewrite /modv eprodv_addl.
apply: (subsetv_trans (addvS Hm1 (subsetv_refl _))).
exact: (addvS (subsetv_refl _) Hm2).
Qed.

Lemma modv_cap : forall ms1 ms2 al , 
  modv ms1 al -> modv ms2 al -> modv (ms1:&: ms2)%VS al.
Proof.
move=> ms1 ms2 al Hm1 Hm2.
by rewrite /modv sub_capv; apply/andP; split;
  [apply: subsetv_trans Hm1 | apply: subsetv_trans Hm2]; 
   apply: eprodv_monol; rewrite (capvSr,capvSl).
Qed.

Definition irreducible ms al := 
  [/\ modv ms al, ms != 0%:VS &
    forall ms1, modv ms1 al -> (ms1 <= ms)%VS -> ms != 0%:VS -> ms1 = ms].

Definition completely_reducible ms al := 
  forall ms1, modv ms1 al -> (ms1 <= ms)%VS -> 
    exists ms2, 
    [/\ modv ms2 al, (ms1 :&: ms2 = 0%:VS)%VS & (ms1 + ms2)%VS = ms].

Lemma completely_reducible0 : forall al, completely_reducible 0%:VS al.
Proof.
move=> al ms1 Hms1; rewrite subsetv0; move/eqP->.
by exists 0%:VS; split; [exact: mod0v | exact: cap0v | exact: sum0v].
Qed.

End AModuleDef.

Notation "a :* b" := (rmul a b): ring_scope.
Notation "A :* B" := (eprodv A B) : vspace_scope.

Module LApp.

Section LinearAppStruct.

(* Endomorphisms over V have an algebra structure as soon as dim V != 0 *)
Variable (R : comRingType) (V: vectType R).
Hypothesis dim_nz: (vdim V != 0)%N.

Canonical Structure algType := LApp.algType dim_nz.

Canonical Structure algFType := Eval hnf in AlgFType R (linearMixin V V).
 
End LinearAppStruct.

End LApp.

Section HomMorphism.

Variable (K: fieldType) (A: algFType K) (M1 M2: amoduleType A).

Implicit Types ms : {vspace M1}.
Implicit Types f : 'Hom(M1, M2).
Implicit Types al : {algebra A}.

Definition modf f ms al :=
       all (fun p => f (p.1 :* p.2) == f p.1 :* p.2) 
               (allpairs (fun x y => (x,y)) (vbasis ms) (vbasis al)).

Lemma modfP : forall f ms al, 
  reflect (forall x v, v \in ms -> x \in al ->  f (v :* x) = f v :* x) 
          (modf f ms al).
Proof.
move=> f ms al; apply: (iffP idP)=> H; last first.
  apply/allP=> [] [v x]; case/allpairsP=> [[x1 x2] [I1 I2 ->]].
  by apply/eqP; apply: H; apply: memv_basis.
move=> x v Hv Hx; rewrite (coord_basis Hv) (coord_basis Hx).
rewrite !linear_sum; apply: eq_big=> //= i _.
rewrite !linearZ /=; congr (_ *: _).
rewrite -!rmul_sum linear_sum; apply: eq_big=> //= j _.
rewrite rmulZ !linearZ /= rmulZ; congr (_ *: _).
set x1 := _`_ _; set y1 := _ `_ _.
case: f H => f /=; move/allP; move/(_ (x1,y1))=> HH.
apply/eqP; apply: HH; apply/allpairsP; exists (x1, y1).
by rewrite !mem_nth /=.
Qed.

Lemma modf_zero : forall ms al, modf 0 ms al.
Proof. by move=> ms al; apply/allP=> i _; rewrite !lappE rmul0. Qed.

Lemma modf_add : forall f1 f2 ms al, 
  modf f1 ms al -> modf f2 ms al -> modf (f1 + f2) ms al.
Proof.
move=> f1 f2 ms al Hm1 Hm2; apply/allP=> [] [v x].
case/allpairsP=> [[x1 x2] [I1 I2 ->]]; rewrite !lappE rmulD.
move/modfP: Hm1->; try apply: memv_basis=>//.
by move/modfP: Hm2->; try apply: memv_basis.
Qed.

Lemma modf_scale : forall k f ms al, modf f ms al -> modf (k *: f) ms al.
Proof.
move=> k f ms al Hm; apply/allP=>  [] [v x].
case/allpairsP=> [[x1 x2] [I1 I2 ->]]; rewrite !lappE rmulZ.
by move/modfP: Hm->; try apply: memv_basis.
Qed.

Lemma modv_ker : forall f ms al, 
  modv ms al -> modf f ms al -> modv (ms :&: lker f)%VS al.
Proof.
move=> f ms al Hmd Hmf; apply/eprodvP=> x v.
rewrite memv_cap !memv_ker.
case/andP=> Hx Hf Hv.
rewrite memv_cap (memv_mod_mul Hmd) // memv_ker.
by move/modfP: Hmf=> ->; rewrite // (eqP Hf) rmul0 eqxx.
Qed.

Lemma modv_img : forall f ms al, 
  modv ms al -> modf f ms al -> modv (f @: ms)%VS al.
Proof.
move=> f ms al Hmv Hmf; apply/eprodvP=> v x.
case/memv_imgP=> u [Hu ->] Hx.
move/modfP: Hmf<-=> //.
apply: memv_img.
by apply: (memv_mod_mul Hmv).
Qed.

End HomMorphism.

Section ModuleRepresentation.

Variable (F: fieldType) (gT: finGroupType) 
         (G: {group gT}) (M: amoduleType (galg F gT)).
Hypothesis CG: ([char F]^'.-group G)%g.
Implicit Types ms : {vspace M}.

Let FG := gaspace F G.
Local Notation " g %:FG " := (injG _ g).

Lemma Maschke : forall ms, modv ms FG -> completely_reducible ms FG.
Proof.
move=> ms Hmv ms1 Hms1 Hsub; rewrite /completely_reducible.
pose act g : 'End(M) := rmorph M (g%:FG).
have actE: forall g v, act g v  = v :* g%:FG by done.
pose f: 'End(M) :=  (#|G|%:R^-1 \*: 
        (\sum_(i \in G) (act (i^-1)%g \o projv ms1 \o (act i))%VS)%R)%VS.
have Cf: forall v x, x \in FG -> f (v :* x) = f v :* x.
  move=> v x; case/memv_sumP=> g_ [Hg_ ->].
  rewrite !linear_sum; apply: eq_big => //= i Hi.
  move: (Hg_ _ Hi); case/injvP=> k ->.
  rewrite !linearZ /=; congr (_ *: _).
  rewrite /f /= !lappE rmulZ; congr (_ *: _).
  rewrite -rmul_sum (reindex (fun g => (i^-1 * g)%g)); last first.
    by exists (fun g => (i * g)%g)=> h; rewrite mulgA (mulVg, mulgV) mul1g.
  apply: eq_big=> g; first by rewrite groupMl // groupV.
  rewrite !lappE /= !lappE /= !actE -rmulA=> Hig.
  have Hg: g \in G by rewrite -[g]mul1g -[1%g](mulgV i) -mulgA groupM.
  by rewrite -injGM // mulgA mulgV mul1g invMg invgK !injGM
             ?groupV // rmulA.
have Himf: forall v, v \in ms1 -> f v = v.
  move=> v Hv.
  rewrite /f !lappE (eq_bigr (fun x => v)); last move=> i Hi.
    by rewrite sumr_const -scaler_nat scalerA mulVf // ?scale1r // -?charf'_nat.
  rewrite !lappE /= !lappE /= projv_id !actE; last first.
    by rewrite (memv_mod_mul Hms1) // /in_mem /= /gvspace (bigD1 i) //=  addvSl.
  by rewrite -rmulA -injGM // ?groupV // mulgV rmul1.
have If: limg f = ms1.
  apply: subsetv_anti; apply/andP; split; last first.
    by apply/subsetvP=> v Hv; rewrite limgE -(Himf _ Hv) memv_img // memvf.
  rewrite limgE; apply/subsetvP=> i; case/memv_imgP=> x [_ ->].
  rewrite !lappE memvZl // memv_sum=> // j Hj.
  rewrite lappE /= lappE (memv_mod_mul Hms1) //; first by exact: memv_proj.
  by rewrite  /in_mem /= /gaspace /gvspace (bigD1 (j^-1)%g) ?addvSl // groupV.
exists (ms :&: lker f)%VS; split.
  - apply: modv_ker=> //; apply/modfP=> *; exact: Cf.
  apply/eqP; rewrite -subsetv0; apply/subsetvP=> v; rewrite memv0.
  rewrite !memv_cap; case/andP=> Hv1; case/andP=> Hv2 Hv3.
  by move: Hv3; rewrite memv_ker  Himf.
apply: subsetv_anti; rewrite  addv_sub Hsub capvSl.
apply/subsetvP=> v Hv.
have->: v = f v + (v - f v) by rewrite addrC -addrA addNr addr0.
apply: addv_mem; first by rewrite -If limgE memv_img // memvf.
rewrite memv_cap; apply/andP; split.
  apply: memv_sub=> //; apply: subsetv_trans Hsub.
  by rewrite -If limgE; apply: memv_img; exact: memvf.
rewrite memv_ker linear_sub /= (Himf (f v)) ?subrr // /in_mem /= -If limgE.
by apply: memv_img; exact: memvf. 
Qed.

End ModuleRepresentation.

Export AModuleType.Exports.